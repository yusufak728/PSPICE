*Yusuf Ahmed Khan 20ELB084

Vcc 3 0 DC 15V
Rc 3 2 1K
Rb 4 1 10K
R1 3 4 12K
R2 4 0 1K
C1 4 5 10UF
VIN 5 0 SIN (0 10M 1K)
Q1 2 1 0 Q2N2222
.model Q2N2222	NPN(Is=14.34f Xti=3 Eg=1.11 Vaf=74.03 Bf=255.9 Ne=1.307
+		Ise=14.34f Ikf=.2847 Xtb=1.5 Br=6.092 Nc=2 Isc=0 Ikr=0 Rc=1
+		Cjc=7.306p Mjc=.3416 Vjc=.75 Fc=.5 Cje=22.01p Mje=.377 Vje=.75
+		Tr=46.91n Tf=411.1p Itf=.6 Vtf=1.7 Xtf=3 Rb=10)
.TRAN 0.1U 5M
.PROBE
.END
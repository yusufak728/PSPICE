*Yusuf Ahmed Khan 20ELB084

Vcc 3 0 DC 15V
Rc 3 2 15K
Rb 4 1 10K
Vbb 4 0 DC 7V
Qt 2 1 0 Q2N2222
.model Q2N2222 npn()
.PROBE
.END
* Yusuf Ahmed Khan
*VIN 6 1 SIN(0 1 1K)
*VDC 1 0 0
*R1 6 2 1k
*R2 2 5 10K
*VP 3 1 15
*VN 4 1 -15
*X1 1 2 3 4 5 UA741

V+ 3 0 5
V- 4 0 -5
X 1 2 3 4 5 UA741

* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt uA741    1 2 3 4 5
*
c1   11 12 8.661E-12
c2    6  7 30.00E-12
dc    5 53 dy
de   54  5 dy
dlp  90 91 dx
dln  92 90 dx
dp    4  3 dx
egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
fb    7 99 poly(5) vb vc ve vlp vln 0 10.61E6 -1E3 1E3 10E6 -10E6
ga    6  0 11 12 188.5E-6
gcm   0  6 10 99 5.961E-9
iee  10  4 dc 15.16E-6
hlim 90  0 vlim 1K
q1   11  2 13 qx
q2   12  1 14 qx
r2    6  9 100.0E3
rc1   3 11 5.305E3
rc2   3 12 5.305E3
re1  13 10 1.836E3
re2  14 10 1.836E3
ree  10 99 13.19E6
ro1   8  5 50
ro2   7 99 100
rp    3  4 18.16E3
vb    9  0 dc 0
vc    3 53 dc 1
ve   54  4 dc 1
vlim  7  8 dc 0
vlp  91  0 dc 40
vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
RG 2 0 10K
RF 5 2 200K
C1 5 6 0.01U
R1 6 1 1.769K
C2 1 0 0.01U
R2 1 0 1.769K
*.FOUR 1K V(5)
.TRAN 0.1MS 2MS
.PROBE
.END




--------------------------------------------------------------------------
